MACRO FD
  ORIGIN 0 0 ;
  FOREIGN FD 0 0 ;
  SIZE 5.16 BY 60.48 ;
  PIN VOUT
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 3.7 2.8 4.9 3.08 ;
      LAYER M2 ;
        RECT 3.7 12.04 4.9 12.32 ;
      LAYER M2 ;
        RECT 3.71 2.8 4.03 3.08 ;
      LAYER M3 ;
        RECT 3.73 2.94 4.01 12.18 ;
      LAYER M2 ;
        RECT 3.71 12.04 4.03 12.32 ;
      LAYER M2 ;
        RECT 1.98 23.38 3.18 23.66 ;
      LAYER M2 ;
        RECT 1.98 21.7 3.18 21.98 ;
      LAYER M2 ;
        RECT 2.42 23.38 2.74 23.66 ;
      LAYER M3 ;
        RECT 2.44 21.84 2.72 23.52 ;
      LAYER M2 ;
        RECT 2.42 21.7 2.74 21.98 ;
      LAYER M2 ;
        RECT 3.44 12.04 3.87 12.32 ;
      LAYER M1 ;
        RECT 3.315 12.18 3.565 21.84 ;
      LAYER M2 ;
        RECT 3.01 21.7 3.44 21.98 ;
    END
  END VOUT
  PIN CLKB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 1.55 27.16 2.75 27.44 ;
      LAYER M2 ;
        RECT 1.55 42.28 2.75 42.56 ;
      LAYER M2 ;
        RECT 1.29 27.16 1.72 27.44 ;
      LAYER M1 ;
        RECT 1.165 27.3 1.415 42.42 ;
      LAYER M2 ;
        RECT 1.29 42.28 1.72 42.56 ;
    END
  END CLKB
  PIN CLK
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 1.55 17.92 2.75 18.2 ;
      LAYER M2 ;
        RECT 1.55 33.04 2.75 33.32 ;
      LAYER M2 ;
        RECT 1.56 17.92 1.88 18.2 ;
      LAYER M1 ;
        RECT 1.595 18.06 1.845 33.18 ;
      LAYER M2 ;
        RECT 1.56 33.04 1.88 33.32 ;
    END
  END CLK
  OBS 
  LAYER M3 ;
        RECT 3.3 0.68 3.58 6.88 ;
  LAYER M3 ;
        RECT 1.58 0.68 1.86 6.88 ;
  LAYER M3 ;
        RECT 3.3 3.595 3.58 3.965 ;
  LAYER M2 ;
        RECT 1.72 3.64 3.44 3.92 ;
  LAYER M3 ;
        RECT 1.58 3.595 1.86 3.965 ;
  LAYER M3 ;
        RECT 2.87 46.04 3.15 52.24 ;
  LAYER M2 ;
        RECT 1.55 29.26 2.75 29.54 ;
  LAYER M2 ;
        RECT 1.55 30.94 2.75 31.22 ;
  LAYER M3 ;
        RECT 3.3 6.72 3.58 7.56 ;
  LAYER M4 ;
        RECT 3.01 7.16 3.44 7.96 ;
  LAYER M3 ;
        RECT 2.87 7.56 3.15 46.2 ;
  LAYER M3 ;
        RECT 2.87 29.215 3.15 29.585 ;
  LAYER M2 ;
        RECT 2.58 29.26 3.01 29.54 ;
  LAYER M3 ;
        RECT 2.87 30.895 3.15 31.265 ;
  LAYER M2 ;
        RECT 2.58 30.94 3.01 31.22 ;
  LAYER M3 ;
        RECT 2.87 7.375 3.15 7.745 ;
  LAYER M4 ;
        RECT 2.845 7.16 3.175 7.96 ;
  LAYER M3 ;
        RECT 3.3 7.375 3.58 7.745 ;
  LAYER M4 ;
        RECT 3.275 7.16 3.605 7.96 ;
  LAYER M3 ;
        RECT 2.87 7.375 3.15 7.745 ;
  LAYER M4 ;
        RECT 2.845 7.16 3.175 7.96 ;
  LAYER M3 ;
        RECT 3.3 7.375 3.58 7.745 ;
  LAYER M4 ;
        RECT 3.275 7.16 3.605 7.96 ;
  LAYER M2 ;
        RECT 2.85 29.26 3.17 29.54 ;
  LAYER M3 ;
        RECT 2.87 29.24 3.15 29.56 ;
  LAYER M3 ;
        RECT 2.87 7.375 3.15 7.745 ;
  LAYER M4 ;
        RECT 2.845 7.16 3.175 7.96 ;
  LAYER M3 ;
        RECT 3.3 7.375 3.58 7.745 ;
  LAYER M4 ;
        RECT 3.275 7.16 3.605 7.96 ;
  LAYER M2 ;
        RECT 2.85 29.26 3.17 29.54 ;
  LAYER M3 ;
        RECT 2.87 29.24 3.15 29.56 ;
  LAYER M3 ;
        RECT 2.87 7.375 3.15 7.745 ;
  LAYER M4 ;
        RECT 2.845 7.16 3.175 7.96 ;
  LAYER M3 ;
        RECT 3.3 7.375 3.58 7.745 ;
  LAYER M4 ;
        RECT 3.275 7.16 3.605 7.96 ;
  LAYER M2 ;
        RECT 2.85 29.26 3.17 29.54 ;
  LAYER M3 ;
        RECT 2.87 29.24 3.15 29.56 ;
  LAYER M2 ;
        RECT 2.85 30.94 3.17 31.22 ;
  LAYER M3 ;
        RECT 2.87 30.92 3.15 31.24 ;
  LAYER M3 ;
        RECT 2.87 7.375 3.15 7.745 ;
  LAYER M4 ;
        RECT 2.845 7.16 3.175 7.96 ;
  LAYER M3 ;
        RECT 3.3 7.375 3.58 7.745 ;
  LAYER M4 ;
        RECT 3.275 7.16 3.605 7.96 ;
  LAYER M2 ;
        RECT 2.85 29.26 3.17 29.54 ;
  LAYER M3 ;
        RECT 2.87 29.24 3.15 29.56 ;
  LAYER M2 ;
        RECT 2.85 30.94 3.17 31.22 ;
  LAYER M3 ;
        RECT 2.87 30.92 3.15 31.24 ;
  LAYER M3 ;
        RECT 2.87 7.375 3.15 7.745 ;
  LAYER M4 ;
        RECT 2.845 7.16 3.175 7.96 ;
  LAYER M3 ;
        RECT 3.3 7.375 3.58 7.745 ;
  LAYER M4 ;
        RECT 3.275 7.16 3.605 7.96 ;
  LAYER M3 ;
        RECT 3.3 8.24 3.58 14.44 ;
  LAYER M3 ;
        RECT 1.58 8.24 1.86 14.44 ;
  LAYER M3 ;
        RECT 3.3 11.155 3.58 11.525 ;
  LAYER M2 ;
        RECT 1.72 11.2 3.44 11.48 ;
  LAYER M3 ;
        RECT 1.58 11.155 1.86 11.525 ;
  LAYER M3 ;
        RECT 2.87 53.6 3.15 59.8 ;
  LAYER M2 ;
        RECT 1.55 15.82 2.75 16.1 ;
  LAYER M2 ;
        RECT 1.55 44.38 2.75 44.66 ;
  LAYER M3 ;
        RECT 3.3 14.28 3.58 52.92 ;
  LAYER M2 ;
        RECT 3.01 52.78 3.44 53.06 ;
  LAYER M3 ;
        RECT 2.87 52.92 3.15 53.76 ;
  LAYER M3 ;
        RECT 3.3 15.775 3.58 16.145 ;
  LAYER M2 ;
        RECT 2.58 15.82 3.44 16.1 ;
  LAYER M3 ;
        RECT 3.3 44.335 3.58 44.705 ;
  LAYER M2 ;
        RECT 2.58 44.38 3.44 44.66 ;
  LAYER M2 ;
        RECT 2.85 52.78 3.17 53.06 ;
  LAYER M3 ;
        RECT 2.87 52.76 3.15 53.08 ;
  LAYER M2 ;
        RECT 3.28 52.78 3.6 53.06 ;
  LAYER M3 ;
        RECT 3.3 52.76 3.58 53.08 ;
  LAYER M2 ;
        RECT 2.85 52.78 3.17 53.06 ;
  LAYER M3 ;
        RECT 2.87 52.76 3.15 53.08 ;
  LAYER M2 ;
        RECT 3.28 52.78 3.6 53.06 ;
  LAYER M3 ;
        RECT 3.3 52.76 3.58 53.08 ;
  LAYER M2 ;
        RECT 2.85 52.78 3.17 53.06 ;
  LAYER M3 ;
        RECT 2.87 52.76 3.15 53.08 ;
  LAYER M2 ;
        RECT 3.28 15.82 3.6 16.1 ;
  LAYER M3 ;
        RECT 3.3 15.8 3.58 16.12 ;
  LAYER M2 ;
        RECT 3.28 52.78 3.6 53.06 ;
  LAYER M3 ;
        RECT 3.3 52.76 3.58 53.08 ;
  LAYER M2 ;
        RECT 2.85 52.78 3.17 53.06 ;
  LAYER M3 ;
        RECT 2.87 52.76 3.15 53.08 ;
  LAYER M2 ;
        RECT 3.28 15.82 3.6 16.1 ;
  LAYER M3 ;
        RECT 3.3 15.8 3.58 16.12 ;
  LAYER M2 ;
        RECT 3.28 52.78 3.6 53.06 ;
  LAYER M3 ;
        RECT 3.3 52.76 3.58 53.08 ;
  LAYER M2 ;
        RECT 2.85 52.78 3.17 53.06 ;
  LAYER M3 ;
        RECT 2.87 52.76 3.15 53.08 ;
  LAYER M2 ;
        RECT 3.28 15.82 3.6 16.1 ;
  LAYER M3 ;
        RECT 3.3 15.8 3.58 16.12 ;
  LAYER M2 ;
        RECT 3.28 44.38 3.6 44.66 ;
  LAYER M3 ;
        RECT 3.3 44.36 3.58 44.68 ;
  LAYER M2 ;
        RECT 3.28 52.78 3.6 53.06 ;
  LAYER M3 ;
        RECT 3.3 52.76 3.58 53.08 ;
  LAYER M2 ;
        RECT 2.85 52.78 3.17 53.06 ;
  LAYER M3 ;
        RECT 2.87 52.76 3.15 53.08 ;
  LAYER M2 ;
        RECT 3.28 15.82 3.6 16.1 ;
  LAYER M3 ;
        RECT 3.3 15.8 3.58 16.12 ;
  LAYER M2 ;
        RECT 3.28 44.38 3.6 44.66 ;
  LAYER M3 ;
        RECT 3.3 44.36 3.58 44.68 ;
  LAYER M2 ;
        RECT 3.28 52.78 3.6 53.06 ;
  LAYER M3 ;
        RECT 3.3 52.76 3.58 53.08 ;
  LAYER M2 ;
        RECT 0.26 7 1.46 7.28 ;
  LAYER M2 ;
        RECT 0.26 7.84 1.46 8.12 ;
  LAYER M2 ;
        RECT 0.7 7 1.02 7.28 ;
  LAYER M3 ;
        RECT 0.72 7.14 1 7.98 ;
  LAYER M2 ;
        RECT 0.7 7.84 1.02 8.12 ;
  LAYER M2 ;
        RECT 1.55 37.24 2.75 37.52 ;
  LAYER M2 ;
        RECT 1.55 38.08 2.75 38.36 ;
  LAYER M2 ;
        RECT 1.99 37.24 2.31 37.52 ;
  LAYER M3 ;
        RECT 2.01 37.38 2.29 38.22 ;
  LAYER M2 ;
        RECT 1.99 38.08 2.31 38.36 ;
  LAYER M2 ;
        RECT 1.13 7.84 1.45 8.12 ;
  LAYER M3 ;
        RECT 1.15 7.98 1.43 37.38 ;
  LAYER M2 ;
        RECT 1.29 37.24 1.72 37.52 ;
  LAYER M2 ;
        RECT 1.13 7.84 1.45 8.12 ;
  LAYER M3 ;
        RECT 1.15 7.82 1.43 8.14 ;
  LAYER M2 ;
        RECT 1.13 37.24 1.45 37.52 ;
  LAYER M3 ;
        RECT 1.15 37.22 1.43 37.54 ;
  LAYER M2 ;
        RECT 1.13 7.84 1.45 8.12 ;
  LAYER M3 ;
        RECT 1.15 7.82 1.43 8.14 ;
  LAYER M2 ;
        RECT 1.13 37.24 1.45 37.52 ;
  LAYER M3 ;
        RECT 1.15 37.22 1.43 37.54 ;
  LAYER M2 ;
        RECT 1.55 48.16 2.75 48.44 ;
  LAYER M2 ;
        RECT 1.55 57.4 2.75 57.68 ;
  LAYER M2 ;
        RECT 1.56 48.16 1.88 48.44 ;
  LAYER M1 ;
        RECT 1.595 48.3 1.845 57.54 ;
  LAYER M2 ;
        RECT 1.56 57.4 1.88 57.68 ;
  LAYER M2 ;
        RECT 1.98 36.82 3.18 37.1 ;
  LAYER M2 ;
        RECT 1.98 38.5 3.18 38.78 ;
  LAYER M2 ;
        RECT 2.42 36.82 2.74 37.1 ;
  LAYER M3 ;
        RECT 2.44 36.96 2.72 38.64 ;
  LAYER M2 ;
        RECT 2.42 38.5 2.74 38.78 ;
  LAYER M1 ;
        RECT 1.595 38.64 1.845 48.3 ;
  LAYER M2 ;
        RECT 1.72 38.5 2.15 38.78 ;
  LAYER M1 ;
        RECT 1.595 38.555 1.845 38.725 ;
  LAYER M2 ;
        RECT 1.55 38.5 1.89 38.78 ;
  LAYER M1 ;
        RECT 1.595 38.555 1.845 38.725 ;
  LAYER M2 ;
        RECT 1.55 38.5 1.89 38.78 ;
  LAYER M2 ;
        RECT 1.55 52.36 2.75 52.64 ;
  LAYER M2 ;
        RECT 1.55 53.2 2.75 53.48 ;
  LAYER M2 ;
        RECT 1.99 52.36 2.31 52.64 ;
  LAYER M3 ;
        RECT 2.01 52.5 2.29 53.34 ;
  LAYER M2 ;
        RECT 1.99 53.2 2.31 53.48 ;
  LAYER M2 ;
        RECT 1.55 22.96 2.75 23.24 ;
  LAYER M2 ;
        RECT 1.55 22.12 2.75 22.4 ;
  LAYER M2 ;
        RECT 1.99 22.96 2.31 23.24 ;
  LAYER M3 ;
        RECT 2.01 22.26 2.29 23.1 ;
  LAYER M2 ;
        RECT 1.99 22.12 2.31 22.4 ;
  LAYER M2 ;
        RECT 1.56 52.36 1.88 52.64 ;
  LAYER M3 ;
        RECT 1.58 23.1 1.86 52.5 ;
  LAYER M2 ;
        RECT 1.56 22.96 1.88 23.24 ;
  LAYER M2 ;
        RECT 1.56 22.96 1.88 23.24 ;
  LAYER M3 ;
        RECT 1.58 22.94 1.86 23.26 ;
  LAYER M2 ;
        RECT 1.56 52.36 1.88 52.64 ;
  LAYER M3 ;
        RECT 1.58 52.34 1.86 52.66 ;
  LAYER M2 ;
        RECT 1.56 22.96 1.88 23.24 ;
  LAYER M3 ;
        RECT 1.58 22.94 1.86 23.26 ;
  LAYER M2 ;
        RECT 1.56 52.36 1.88 52.64 ;
  LAYER M3 ;
        RECT 1.58 52.34 1.86 52.66 ;
  LAYER M2 ;
        RECT 3.7 7 4.9 7.28 ;
  LAYER M2 ;
        RECT 3.7 7.84 4.9 8.12 ;
  LAYER M2 ;
        RECT 4.14 7 4.46 7.28 ;
  LAYER M3 ;
        RECT 4.16 7.14 4.44 7.98 ;
  LAYER M2 ;
        RECT 4.14 7.84 4.46 8.12 ;
  LAYER M2 ;
        RECT 0.26 2.8 1.46 3.08 ;
  LAYER M2 ;
        RECT 0.26 12.04 1.46 12.32 ;
  LAYER M2 ;
        RECT 0.27 2.8 0.59 3.08 ;
  LAYER M1 ;
        RECT 0.305 2.94 0.555 12.18 ;
  LAYER M2 ;
        RECT 0.27 12.04 0.59 12.32 ;
  LAYER M3 ;
        RECT 4.16 7.375 4.44 7.745 ;
  LAYER M2 ;
        RECT 0.43 7.42 4.3 7.7 ;
  LAYER M1 ;
        RECT 0.305 7.475 0.555 7.645 ;
  LAYER M1 ;
        RECT 0.305 7.475 0.555 7.645 ;
  LAYER M2 ;
        RECT 0.26 7.42 0.6 7.7 ;
  LAYER M2 ;
        RECT 4.14 7.42 4.46 7.7 ;
  LAYER M3 ;
        RECT 4.16 7.4 4.44 7.72 ;
  LAYER M1 ;
        RECT 0.305 7.475 0.555 7.645 ;
  LAYER M2 ;
        RECT 0.26 7.42 0.6 7.7 ;
  LAYER M2 ;
        RECT 4.14 7.42 4.46 7.7 ;
  LAYER M3 ;
        RECT 4.16 7.4 4.44 7.72 ;
  LAYER M1 ;
        RECT 3.745 3.695 3.995 7.225 ;
  LAYER M1 ;
        RECT 3.745 2.435 3.995 3.445 ;
  LAYER M1 ;
        RECT 3.745 0.335 3.995 1.345 ;
  LAYER M1 ;
        RECT 4.175 3.695 4.425 7.225 ;
  LAYER M1 ;
        RECT 3.315 3.695 3.565 7.225 ;
  LAYER M2 ;
        RECT 3.27 0.7 4.47 0.98 ;
  LAYER M2 ;
        RECT 3.27 6.58 4.47 6.86 ;
  LAYER M2 ;
        RECT 3.7 7 4.9 7.28 ;
  LAYER M2 ;
        RECT 3.7 2.8 4.9 3.08 ;
  LAYER M3 ;
        RECT 3.3 0.68 3.58 6.88 ;
  LAYER M1 ;
        RECT 3.745 7.895 3.995 11.425 ;
  LAYER M1 ;
        RECT 3.745 11.675 3.995 12.685 ;
  LAYER M1 ;
        RECT 3.745 13.775 3.995 14.785 ;
  LAYER M1 ;
        RECT 4.175 7.895 4.425 11.425 ;
  LAYER M1 ;
        RECT 3.315 7.895 3.565 11.425 ;
  LAYER M2 ;
        RECT 3.27 14.14 4.47 14.42 ;
  LAYER M2 ;
        RECT 3.27 8.26 4.47 8.54 ;
  LAYER M2 ;
        RECT 3.7 7.84 4.9 8.12 ;
  LAYER M2 ;
        RECT 3.7 12.04 4.9 12.32 ;
  LAYER M3 ;
        RECT 3.3 8.24 3.58 14.44 ;
  LAYER M1 ;
        RECT 1.165 3.695 1.415 7.225 ;
  LAYER M1 ;
        RECT 1.165 2.435 1.415 3.445 ;
  LAYER M1 ;
        RECT 1.165 0.335 1.415 1.345 ;
  LAYER M1 ;
        RECT 0.735 3.695 0.985 7.225 ;
  LAYER M1 ;
        RECT 1.595 3.695 1.845 7.225 ;
  LAYER M2 ;
        RECT 0.69 0.7 1.89 0.98 ;
  LAYER M2 ;
        RECT 0.69 6.58 1.89 6.86 ;
  LAYER M2 ;
        RECT 0.26 7 1.46 7.28 ;
  LAYER M2 ;
        RECT 0.26 2.8 1.46 3.08 ;
  LAYER M3 ;
        RECT 1.58 0.68 1.86 6.88 ;
  LAYER M1 ;
        RECT 1.165 7.895 1.415 11.425 ;
  LAYER M1 ;
        RECT 1.165 11.675 1.415 12.685 ;
  LAYER M1 ;
        RECT 1.165 13.775 1.415 14.785 ;
  LAYER M1 ;
        RECT 0.735 7.895 0.985 11.425 ;
  LAYER M1 ;
        RECT 1.595 7.895 1.845 11.425 ;
  LAYER M2 ;
        RECT 0.69 14.14 1.89 14.42 ;
  LAYER M2 ;
        RECT 0.69 8.26 1.89 8.54 ;
  LAYER M2 ;
        RECT 0.26 7.84 1.46 8.12 ;
  LAYER M2 ;
        RECT 0.26 12.04 1.46 12.32 ;
  LAYER M3 ;
        RECT 1.58 8.24 1.86 14.44 ;
  LAYER M1 ;
        RECT 2.455 49.055 2.705 52.585 ;
  LAYER M1 ;
        RECT 2.455 47.795 2.705 48.805 ;
  LAYER M1 ;
        RECT 2.455 45.695 2.705 46.705 ;
  LAYER M1 ;
        RECT 2.025 49.055 2.275 52.585 ;
  LAYER M1 ;
        RECT 2.885 49.055 3.135 52.585 ;
  LAYER M2 ;
        RECT 1.98 46.06 3.18 46.34 ;
  LAYER M2 ;
        RECT 1.98 51.94 3.18 52.22 ;
  LAYER M2 ;
        RECT 1.55 52.36 2.75 52.64 ;
  LAYER M2 ;
        RECT 1.55 48.16 2.75 48.44 ;
  LAYER M3 ;
        RECT 2.87 46.04 3.15 52.24 ;
  LAYER M1 ;
        RECT 2.455 53.255 2.705 56.785 ;
  LAYER M1 ;
        RECT 2.455 57.035 2.705 58.045 ;
  LAYER M1 ;
        RECT 2.455 59.135 2.705 60.145 ;
  LAYER M1 ;
        RECT 2.025 53.255 2.275 56.785 ;
  LAYER M1 ;
        RECT 2.885 53.255 3.135 56.785 ;
  LAYER M2 ;
        RECT 1.98 59.5 3.18 59.78 ;
  LAYER M2 ;
        RECT 1.98 53.62 3.18 53.9 ;
  LAYER M2 ;
        RECT 1.55 53.2 2.75 53.48 ;
  LAYER M2 ;
        RECT 1.55 57.4 2.75 57.68 ;
  LAYER M3 ;
        RECT 2.87 53.6 3.15 59.8 ;
  LAYER M1 ;
        RECT 2.455 23.015 2.705 26.545 ;
  LAYER M1 ;
        RECT 2.455 26.795 2.705 27.805 ;
  LAYER M1 ;
        RECT 2.455 28.895 2.705 29.905 ;
  LAYER M1 ;
        RECT 2.025 23.015 2.275 26.545 ;
  LAYER M1 ;
        RECT 2.885 23.015 3.135 26.545 ;
  LAYER M2 ;
        RECT 1.55 29.26 2.75 29.54 ;
  LAYER M2 ;
        RECT 1.55 22.96 2.75 23.24 ;
  LAYER M2 ;
        RECT 1.55 27.16 2.75 27.44 ;
  LAYER M2 ;
        RECT 1.98 23.38 3.18 23.66 ;
  LAYER M1 ;
        RECT 2.455 18.815 2.705 22.345 ;
  LAYER M1 ;
        RECT 2.455 17.555 2.705 18.565 ;
  LAYER M1 ;
        RECT 2.455 15.455 2.705 16.465 ;
  LAYER M1 ;
        RECT 2.025 18.815 2.275 22.345 ;
  LAYER M1 ;
        RECT 2.885 18.815 3.135 22.345 ;
  LAYER M2 ;
        RECT 1.55 15.82 2.75 16.1 ;
  LAYER M2 ;
        RECT 1.55 22.12 2.75 22.4 ;
  LAYER M2 ;
        RECT 1.55 17.92 2.75 18.2 ;
  LAYER M2 ;
        RECT 1.98 21.7 3.18 21.98 ;
  LAYER M1 ;
        RECT 2.455 33.935 2.705 37.465 ;
  LAYER M1 ;
        RECT 2.455 32.675 2.705 33.685 ;
  LAYER M1 ;
        RECT 2.455 30.575 2.705 31.585 ;
  LAYER M1 ;
        RECT 2.025 33.935 2.275 37.465 ;
  LAYER M1 ;
        RECT 2.885 33.935 3.135 37.465 ;
  LAYER M2 ;
        RECT 1.55 30.94 2.75 31.22 ;
  LAYER M2 ;
        RECT 1.55 37.24 2.75 37.52 ;
  LAYER M2 ;
        RECT 1.55 33.04 2.75 33.32 ;
  LAYER M2 ;
        RECT 1.98 36.82 3.18 37.1 ;
  LAYER M1 ;
        RECT 2.455 38.135 2.705 41.665 ;
  LAYER M1 ;
        RECT 2.455 41.915 2.705 42.925 ;
  LAYER M1 ;
        RECT 2.455 44.015 2.705 45.025 ;
  LAYER M1 ;
        RECT 2.025 38.135 2.275 41.665 ;
  LAYER M1 ;
        RECT 2.885 38.135 3.135 41.665 ;
  LAYER M2 ;
        RECT 1.55 44.38 2.75 44.66 ;
  LAYER M2 ;
        RECT 1.55 38.08 2.75 38.36 ;
  LAYER M2 ;
        RECT 1.55 42.28 2.75 42.56 ;
  LAYER M2 ;
        RECT 1.98 38.5 3.18 38.78 ;
  END 
END FD

MACRO CP
  ORIGIN 0 0 ;
  FOREIGN CP 0 0 ;
  SIZE 11.18 BY 22.68 ;
  PIN VSS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 7.17 16.22 7.45 22 ;
      LAYER M3 ;
        RECT 1.58 8.24 1.86 14.44 ;
      LAYER M3 ;
        RECT 9.32 8.24 9.6 14.44 ;
      LAYER M3 ;
        RECT 9.32 15.8 9.6 22 ;
      LAYER M3 ;
        RECT 7.17 15.12 7.45 16.38 ;
      LAYER M2 ;
        RECT 1.72 14.98 7.31 15.26 ;
      LAYER M3 ;
        RECT 1.58 14.28 1.86 15.12 ;
      LAYER M3 ;
        RECT 7.17 14.935 7.45 15.305 ;
      LAYER M4 ;
        RECT 7.31 14.72 9.46 15.52 ;
      LAYER M3 ;
        RECT 9.32 14.28 9.6 15.12 ;
      LAYER M3 ;
        RECT 9.32 15.12 9.6 15.96 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 7.17 0.68 7.45 6.46 ;
      LAYER M3 ;
        RECT 1.58 0.68 1.86 6.88 ;
      LAYER M3 ;
        RECT 9.32 0.68 9.6 6.88 ;
      LAYER M3 ;
        RECT 4.16 0.68 4.44 6.88 ;
      LAYER M3 ;
        RECT 7.17 3.595 7.45 3.965 ;
      LAYER M2 ;
        RECT 1.72 3.64 7.31 3.92 ;
      LAYER M3 ;
        RECT 1.58 3.595 1.86 3.965 ;
      LAYER M3 ;
        RECT 7.17 3.595 7.45 3.965 ;
      LAYER M4 ;
        RECT 7.31 3.38 9.46 4.18 ;
      LAYER M3 ;
        RECT 9.32 3.595 9.6 3.965 ;
      LAYER M2 ;
        RECT 4.14 3.64 4.46 3.92 ;
      LAYER M3 ;
        RECT 4.16 3.595 4.44 3.965 ;
    END
  END VDD
  PIN UP
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 0.26 7.84 1.46 8.12 ;
      LAYER M2 ;
        RECT 0.26 7 1.46 7.28 ;
      LAYER M2 ;
        RECT 0.7 7.84 1.02 8.12 ;
      LAYER M3 ;
        RECT 0.72 7.14 1 7.98 ;
      LAYER M2 ;
        RECT 0.7 7 1.02 7.28 ;
      LAYER M2 ;
        RECT 0.26 19.6 1.46 19.88 ;
      LAYER M2 ;
        RECT 0.27 7.84 0.59 8.12 ;
      LAYER M3 ;
        RECT 0.29 7.98 0.57 19.74 ;
      LAYER M2 ;
        RECT 0.27 19.6 0.59 19.88 ;
    END
  END UP
  PIN DN
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 9.72 7.84 10.92 8.12 ;
      LAYER M2 ;
        RECT 9.72 7 10.92 7.28 ;
      LAYER M2 ;
        RECT 10.16 7.84 10.48 8.12 ;
      LAYER M3 ;
        RECT 10.18 7.14 10.46 7.98 ;
      LAYER M2 ;
        RECT 10.16 7 10.48 7.28 ;
      LAYER M2 ;
        RECT 7.14 10.36 8.34 10.64 ;
      LAYER M2 ;
        RECT 9.03 7.84 9.89 8.12 ;
      LAYER M1 ;
        RECT 8.905 7.98 9.155 10.5 ;
      LAYER M2 ;
        RECT 8.17 10.36 9.03 10.64 ;
    END
  END DN
  PIN OUT
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 0.26 15.4 1.46 15.68 ;
      LAYER M2 ;
        RECT 3.7 14.56 4.9 14.84 ;
      LAYER M2 ;
        RECT 1.13 15.4 1.45 15.68 ;
      LAYER M3 ;
        RECT 1.15 15.12 1.43 15.54 ;
      LAYER M4 ;
        RECT 1.29 14.72 2.15 15.52 ;
      LAYER M3 ;
        RECT 2.01 14.7 2.29 15.12 ;
      LAYER M2 ;
        RECT 2.15 14.56 3.87 14.84 ;
    END
  END OUT
  OBS 
  LAYER M3 ;
        RECT 6.31 15.38 6.59 19.9 ;
  LAYER M2 ;
        RECT 6.28 15.82 7.48 16.1 ;
  LAYER M3 ;
        RECT 4.16 15.8 4.44 22 ;
  LAYER M3 ;
        RECT 1.58 15.8 1.86 22 ;
  LAYER M2 ;
        RECT 5.16 15.82 6.45 16.1 ;
  LAYER M1 ;
        RECT 5.035 15.96 5.285 16.38 ;
  LAYER M2 ;
        RECT 4.3 16.24 5.16 16.52 ;
  LAYER M3 ;
        RECT 4.16 16.195 4.44 16.565 ;
  LAYER M3 ;
        RECT 4.16 18.715 4.44 19.085 ;
  LAYER M2 ;
        RECT 1.72 18.76 4.3 19.04 ;
  LAYER M3 ;
        RECT 1.58 18.715 1.86 19.085 ;
  LAYER M1 ;
        RECT 5.035 15.875 5.285 16.045 ;
  LAYER M2 ;
        RECT 4.99 15.82 5.33 16.1 ;
  LAYER M1 ;
        RECT 5.035 16.295 5.285 16.465 ;
  LAYER M2 ;
        RECT 4.99 16.24 5.33 16.52 ;
  LAYER M2 ;
        RECT 4.14 16.24 4.46 16.52 ;
  LAYER M3 ;
        RECT 4.16 16.22 4.44 16.54 ;
  LAYER M1 ;
        RECT 5.035 15.875 5.285 16.045 ;
  LAYER M2 ;
        RECT 4.99 15.82 5.33 16.1 ;
  LAYER M1 ;
        RECT 5.035 16.295 5.285 16.465 ;
  LAYER M2 ;
        RECT 4.99 16.24 5.33 16.52 ;
  LAYER M2 ;
        RECT 4.14 16.24 4.46 16.52 ;
  LAYER M3 ;
        RECT 4.16 16.22 4.44 16.54 ;
  LAYER M1 ;
        RECT 5.035 15.875 5.285 16.045 ;
  LAYER M2 ;
        RECT 4.99 15.82 5.33 16.1 ;
  LAYER M1 ;
        RECT 5.035 16.295 5.285 16.465 ;
  LAYER M2 ;
        RECT 4.99 16.24 5.33 16.52 ;
  LAYER M2 ;
        RECT 1.56 18.76 1.88 19.04 ;
  LAYER M3 ;
        RECT 1.58 18.74 1.86 19.06 ;
  LAYER M2 ;
        RECT 4.14 16.24 4.46 16.52 ;
  LAYER M3 ;
        RECT 4.16 16.22 4.44 16.54 ;
  LAYER M2 ;
        RECT 4.14 18.76 4.46 19.04 ;
  LAYER M3 ;
        RECT 4.16 18.74 4.44 19.06 ;
  LAYER M1 ;
        RECT 5.035 15.875 5.285 16.045 ;
  LAYER M2 ;
        RECT 4.99 15.82 5.33 16.1 ;
  LAYER M1 ;
        RECT 5.035 16.295 5.285 16.465 ;
  LAYER M2 ;
        RECT 4.99 16.24 5.33 16.52 ;
  LAYER M2 ;
        RECT 1.56 18.76 1.88 19.04 ;
  LAYER M3 ;
        RECT 1.58 18.74 1.86 19.06 ;
  LAYER M2 ;
        RECT 4.14 16.24 4.46 16.52 ;
  LAYER M3 ;
        RECT 4.16 16.22 4.44 16.54 ;
  LAYER M2 ;
        RECT 4.14 18.76 4.46 19.04 ;
  LAYER M3 ;
        RECT 4.16 18.74 4.44 19.06 ;
  LAYER M3 ;
        RECT 6.31 2.78 6.59 7.3 ;
  LAYER M2 ;
        RECT 6.28 6.58 7.48 6.86 ;
  LAYER M3 ;
        RECT 5.02 8.24 5.3 14.44 ;
  LAYER M3 ;
        RECT 6.74 8.24 7.02 14.44 ;
  LAYER M2 ;
        RECT 5.16 6.58 6.45 6.86 ;
  LAYER M3 ;
        RECT 5.02 6.72 5.3 8.4 ;
  LAYER M2 ;
        RECT 6.72 6.58 7.04 6.86 ;
  LAYER M3 ;
        RECT 6.74 6.72 7.02 8.4 ;
  LAYER M2 ;
        RECT 5 6.58 5.32 6.86 ;
  LAYER M3 ;
        RECT 5.02 6.56 5.3 6.88 ;
  LAYER M2 ;
        RECT 5 6.58 5.32 6.86 ;
  LAYER M3 ;
        RECT 5.02 6.56 5.3 6.88 ;
  LAYER M2 ;
        RECT 5 6.58 5.32 6.86 ;
  LAYER M3 ;
        RECT 5.02 6.56 5.3 6.88 ;
  LAYER M2 ;
        RECT 6.72 6.58 7.04 6.86 ;
  LAYER M3 ;
        RECT 6.74 6.56 7.02 6.88 ;
  LAYER M2 ;
        RECT 5 6.58 5.32 6.86 ;
  LAYER M3 ;
        RECT 5.02 6.56 5.3 6.88 ;
  LAYER M2 ;
        RECT 6.72 6.58 7.04 6.86 ;
  LAYER M3 ;
        RECT 6.74 6.56 7.02 6.88 ;
  LAYER M2 ;
        RECT 0.26 12.04 1.46 12.32 ;
  LAYER M2 ;
        RECT 0.26 2.8 1.46 3.08 ;
  LAYER M2 ;
        RECT 0.27 12.04 0.59 12.32 ;
  LAYER M1 ;
        RECT 0.305 2.94 0.555 12.18 ;
  LAYER M2 ;
        RECT 0.27 2.8 0.59 3.08 ;
  LAYER M2 ;
        RECT 2.84 19.6 4.04 19.88 ;
  LAYER M2 ;
        RECT 1.29 12.04 2.15 12.32 ;
  LAYER M1 ;
        RECT 2.025 12.18 2.275 19.74 ;
  LAYER M2 ;
        RECT 2.15 19.6 3.01 19.88 ;
  LAYER M1 ;
        RECT 2.025 12.095 2.275 12.265 ;
  LAYER M2 ;
        RECT 1.98 12.04 2.32 12.32 ;
  LAYER M1 ;
        RECT 2.025 19.655 2.275 19.825 ;
  LAYER M2 ;
        RECT 1.98 19.6 2.32 19.88 ;
  LAYER M1 ;
        RECT 2.025 12.095 2.275 12.265 ;
  LAYER M2 ;
        RECT 1.98 12.04 2.32 12.32 ;
  LAYER M1 ;
        RECT 2.025 19.655 2.275 19.825 ;
  LAYER M2 ;
        RECT 1.98 19.6 2.32 19.88 ;
  LAYER M2 ;
        RECT 9.72 12.04 10.92 12.32 ;
  LAYER M2 ;
        RECT 9.72 2.8 10.92 3.08 ;
  LAYER M2 ;
        RECT 9.73 12.04 10.05 12.32 ;
  LAYER M3 ;
        RECT 9.75 2.94 10.03 12.18 ;
  LAYER M2 ;
        RECT 9.73 2.8 10.05 3.08 ;
  LAYER M2 ;
        RECT 3.7 10.36 4.9 10.64 ;
  LAYER M3 ;
        RECT 9.75 9.895 10.03 10.265 ;
  LAYER M2 ;
        RECT 6.45 9.94 9.89 10.22 ;
  LAYER M1 ;
        RECT 6.325 10.08 6.575 10.5 ;
  LAYER M2 ;
        RECT 4.73 10.36 6.45 10.64 ;
  LAYER M1 ;
        RECT 6.325 9.995 6.575 10.165 ;
  LAYER M2 ;
        RECT 6.28 9.94 6.62 10.22 ;
  LAYER M1 ;
        RECT 6.325 10.415 6.575 10.585 ;
  LAYER M2 ;
        RECT 6.28 10.36 6.62 10.64 ;
  LAYER M2 ;
        RECT 9.73 9.94 10.05 10.22 ;
  LAYER M3 ;
        RECT 9.75 9.92 10.03 10.24 ;
  LAYER M1 ;
        RECT 6.325 9.995 6.575 10.165 ;
  LAYER M2 ;
        RECT 6.28 9.94 6.62 10.22 ;
  LAYER M1 ;
        RECT 6.325 10.415 6.575 10.585 ;
  LAYER M2 ;
        RECT 6.28 10.36 6.62 10.64 ;
  LAYER M2 ;
        RECT 9.73 9.94 10.05 10.22 ;
  LAYER M3 ;
        RECT 9.75 9.92 10.03 10.24 ;
  LAYER M3 ;
        RECT 9.75 15.38 10.03 19.9 ;
  LAYER M2 ;
        RECT 7.14 14.56 8.34 14.84 ;
  LAYER M3 ;
        RECT 9.75 16.195 10.03 16.565 ;
  LAYER M2 ;
        RECT 9.03 16.24 9.89 16.52 ;
  LAYER M1 ;
        RECT 8.905 14.7 9.155 16.38 ;
  LAYER M2 ;
        RECT 8.17 14.56 9.03 14.84 ;
  LAYER M1 ;
        RECT 8.905 14.615 9.155 14.785 ;
  LAYER M2 ;
        RECT 8.86 14.56 9.2 14.84 ;
  LAYER M1 ;
        RECT 8.905 16.295 9.155 16.465 ;
  LAYER M2 ;
        RECT 8.86 16.24 9.2 16.52 ;
  LAYER M2 ;
        RECT 9.73 16.24 10.05 16.52 ;
  LAYER M3 ;
        RECT 9.75 16.22 10.03 16.54 ;
  LAYER M1 ;
        RECT 8.905 14.615 9.155 14.785 ;
  LAYER M2 ;
        RECT 8.86 14.56 9.2 14.84 ;
  LAYER M1 ;
        RECT 8.905 16.295 9.155 16.465 ;
  LAYER M2 ;
        RECT 8.86 16.24 9.2 16.52 ;
  LAYER M2 ;
        RECT 9.73 16.24 10.05 16.52 ;
  LAYER M3 ;
        RECT 9.75 16.22 10.03 16.54 ;
  LAYER M3 ;
        RECT 3.73 2.78 4.01 7.3 ;
  LAYER M2 ;
        RECT 2.84 15.4 4.04 15.68 ;
  LAYER M3 ;
        RECT 3.73 7.14 4.01 15.54 ;
  LAYER M2 ;
        RECT 3.71 15.4 4.03 15.68 ;
  LAYER M2 ;
        RECT 3.71 15.4 4.03 15.68 ;
  LAYER M3 ;
        RECT 3.73 15.38 4.01 15.7 ;
  LAYER M2 ;
        RECT 3.71 15.4 4.03 15.68 ;
  LAYER M3 ;
        RECT 3.73 15.38 4.01 15.7 ;
  LAYER M1 ;
        RECT 6.325 15.455 6.575 18.985 ;
  LAYER M1 ;
        RECT 6.325 19.235 6.575 20.245 ;
  LAYER M1 ;
        RECT 6.325 21.335 6.575 22.345 ;
  LAYER M1 ;
        RECT 5.895 15.455 6.145 18.985 ;
  LAYER M1 ;
        RECT 6.755 15.455 7.005 18.985 ;
  LAYER M1 ;
        RECT 7.185 15.455 7.435 18.985 ;
  LAYER M1 ;
        RECT 7.185 19.235 7.435 20.245 ;
  LAYER M1 ;
        RECT 7.185 21.335 7.435 22.345 ;
  LAYER M1 ;
        RECT 7.615 15.455 7.865 18.985 ;
  LAYER M2 ;
        RECT 5.42 15.4 6.62 15.68 ;
  LAYER M2 ;
        RECT 6.28 19.6 7.48 19.88 ;
  LAYER M2 ;
        RECT 5.85 16.24 7.91 16.52 ;
  LAYER M2 ;
        RECT 6.28 21.7 7.48 21.98 ;
  LAYER M3 ;
        RECT 6.31 15.38 6.59 19.9 ;
  LAYER M2 ;
        RECT 6.28 15.82 7.48 16.1 ;
  LAYER M3 ;
        RECT 7.17 16.22 7.45 22 ;
  LAYER M1 ;
        RECT 6.325 3.695 6.575 7.225 ;
  LAYER M1 ;
        RECT 6.325 2.435 6.575 3.445 ;
  LAYER M1 ;
        RECT 6.325 0.335 6.575 1.345 ;
  LAYER M1 ;
        RECT 5.895 3.695 6.145 7.225 ;
  LAYER M1 ;
        RECT 6.755 3.695 7.005 7.225 ;
  LAYER M1 ;
        RECT 7.185 3.695 7.435 7.225 ;
  LAYER M1 ;
        RECT 7.185 2.435 7.435 3.445 ;
  LAYER M1 ;
        RECT 7.185 0.335 7.435 1.345 ;
  LAYER M1 ;
        RECT 7.615 3.695 7.865 7.225 ;
  LAYER M2 ;
        RECT 5.42 7 6.62 7.28 ;
  LAYER M2 ;
        RECT 6.28 2.8 7.48 3.08 ;
  LAYER M2 ;
        RECT 5.85 6.16 7.91 6.44 ;
  LAYER M2 ;
        RECT 6.28 0.7 7.48 0.98 ;
  LAYER M3 ;
        RECT 6.31 2.78 6.59 7.3 ;
  LAYER M2 ;
        RECT 6.28 6.58 7.48 6.86 ;
  LAYER M3 ;
        RECT 7.17 0.68 7.45 6.46 ;
  LAYER M1 ;
        RECT 1.165 7.895 1.415 11.425 ;
  LAYER M1 ;
        RECT 1.165 11.675 1.415 12.685 ;
  LAYER M1 ;
        RECT 1.165 13.775 1.415 14.785 ;
  LAYER M1 ;
        RECT 0.735 7.895 0.985 11.425 ;
  LAYER M1 ;
        RECT 1.595 7.895 1.845 11.425 ;
  LAYER M2 ;
        RECT 0.69 8.26 1.89 8.54 ;
  LAYER M2 ;
        RECT 0.69 14.14 1.89 14.42 ;
  LAYER M2 ;
        RECT 0.26 7.84 1.46 8.12 ;
  LAYER M2 ;
        RECT 0.26 12.04 1.46 12.32 ;
  LAYER M3 ;
        RECT 1.58 8.24 1.86 14.44 ;
  LAYER M1 ;
        RECT 1.165 3.695 1.415 7.225 ;
  LAYER M1 ;
        RECT 1.165 2.435 1.415 3.445 ;
  LAYER M1 ;
        RECT 1.165 0.335 1.415 1.345 ;
  LAYER M1 ;
        RECT 0.735 3.695 0.985 7.225 ;
  LAYER M1 ;
        RECT 1.595 3.695 1.845 7.225 ;
  LAYER M2 ;
        RECT 0.69 6.58 1.89 6.86 ;
  LAYER M2 ;
        RECT 0.69 0.7 1.89 0.98 ;
  LAYER M2 ;
        RECT 0.26 7 1.46 7.28 ;
  LAYER M2 ;
        RECT 0.26 2.8 1.46 3.08 ;
  LAYER M3 ;
        RECT 1.58 0.68 1.86 6.88 ;
  LAYER M1 ;
        RECT 9.765 7.895 10.015 11.425 ;
  LAYER M1 ;
        RECT 9.765 11.675 10.015 12.685 ;
  LAYER M1 ;
        RECT 9.765 13.775 10.015 14.785 ;
  LAYER M1 ;
        RECT 10.195 7.895 10.445 11.425 ;
  LAYER M1 ;
        RECT 9.335 7.895 9.585 11.425 ;
  LAYER M2 ;
        RECT 9.29 8.26 10.49 8.54 ;
  LAYER M2 ;
        RECT 9.29 14.14 10.49 14.42 ;
  LAYER M2 ;
        RECT 9.72 7.84 10.92 8.12 ;
  LAYER M2 ;
        RECT 9.72 12.04 10.92 12.32 ;
  LAYER M3 ;
        RECT 9.32 8.24 9.6 14.44 ;
  LAYER M1 ;
        RECT 9.765 3.695 10.015 7.225 ;
  LAYER M1 ;
        RECT 9.765 2.435 10.015 3.445 ;
  LAYER M1 ;
        RECT 9.765 0.335 10.015 1.345 ;
  LAYER M1 ;
        RECT 10.195 3.695 10.445 7.225 ;
  LAYER M1 ;
        RECT 9.335 3.695 9.585 7.225 ;
  LAYER M2 ;
        RECT 9.29 6.58 10.49 6.86 ;
  LAYER M2 ;
        RECT 9.29 0.7 10.49 0.98 ;
  LAYER M2 ;
        RECT 9.72 7 10.92 7.28 ;
  LAYER M2 ;
        RECT 9.72 2.8 10.92 3.08 ;
  LAYER M3 ;
        RECT 9.32 0.68 9.6 6.88 ;
  LAYER M1 ;
        RECT 9.765 15.455 10.015 18.985 ;
  LAYER M1 ;
        RECT 9.765 19.235 10.015 20.245 ;
  LAYER M1 ;
        RECT 9.765 21.335 10.015 22.345 ;
  LAYER M1 ;
        RECT 10.195 15.455 10.445 18.985 ;
  LAYER M1 ;
        RECT 9.335 15.455 9.585 18.985 ;
  LAYER M2 ;
        RECT 9.72 15.4 10.92 15.68 ;
  LAYER M2 ;
        RECT 9.72 19.6 10.92 19.88 ;
  LAYER M2 ;
        RECT 9.29 15.82 10.49 16.1 ;
  LAYER M2 ;
        RECT 9.29 21.7 10.49 21.98 ;
  LAYER M3 ;
        RECT 9.75 15.38 10.03 19.9 ;
  LAYER M3 ;
        RECT 9.32 15.8 9.6 22 ;
  LAYER M1 ;
        RECT 3.745 3.695 3.995 7.225 ;
  LAYER M1 ;
        RECT 3.745 2.435 3.995 3.445 ;
  LAYER M1 ;
        RECT 3.745 0.335 3.995 1.345 ;
  LAYER M1 ;
        RECT 3.315 3.695 3.565 7.225 ;
  LAYER M1 ;
        RECT 4.175 3.695 4.425 7.225 ;
  LAYER M2 ;
        RECT 2.84 7 4.04 7.28 ;
  LAYER M2 ;
        RECT 2.84 2.8 4.04 3.08 ;
  LAYER M2 ;
        RECT 3.27 6.58 4.47 6.86 ;
  LAYER M2 ;
        RECT 3.27 0.7 4.47 0.98 ;
  LAYER M3 ;
        RECT 3.73 2.78 4.01 7.3 ;
  LAYER M3 ;
        RECT 4.16 0.68 4.44 6.88 ;
  LAYER M1 ;
        RECT 3.745 15.455 3.995 18.985 ;
  LAYER M1 ;
        RECT 3.745 19.235 3.995 20.245 ;
  LAYER M1 ;
        RECT 3.745 21.335 3.995 22.345 ;
  LAYER M1 ;
        RECT 3.315 15.455 3.565 18.985 ;
  LAYER M1 ;
        RECT 4.175 15.455 4.425 18.985 ;
  LAYER M2 ;
        RECT 3.27 15.82 4.47 16.1 ;
  LAYER M2 ;
        RECT 3.27 21.7 4.47 21.98 ;
  LAYER M2 ;
        RECT 2.84 15.4 4.04 15.68 ;
  LAYER M2 ;
        RECT 2.84 19.6 4.04 19.88 ;
  LAYER M3 ;
        RECT 4.16 15.8 4.44 22 ;
  LAYER M1 ;
        RECT 1.165 15.455 1.415 18.985 ;
  LAYER M1 ;
        RECT 1.165 19.235 1.415 20.245 ;
  LAYER M1 ;
        RECT 1.165 21.335 1.415 22.345 ;
  LAYER M1 ;
        RECT 0.735 15.455 0.985 18.985 ;
  LAYER M1 ;
        RECT 1.595 15.455 1.845 18.985 ;
  LAYER M2 ;
        RECT 0.69 15.82 1.89 16.1 ;
  LAYER M2 ;
        RECT 0.69 21.7 1.89 21.98 ;
  LAYER M2 ;
        RECT 0.26 15.4 1.46 15.68 ;
  LAYER M2 ;
        RECT 0.26 19.6 1.46 19.88 ;
  LAYER M3 ;
        RECT 1.58 15.8 1.86 22 ;
  LAYER M1 ;
        RECT 4.605 11.255 4.855 14.785 ;
  LAYER M1 ;
        RECT 4.605 9.995 4.855 11.005 ;
  LAYER M1 ;
        RECT 4.605 7.895 4.855 8.905 ;
  LAYER M1 ;
        RECT 4.175 11.255 4.425 14.785 ;
  LAYER M1 ;
        RECT 5.035 11.255 5.285 14.785 ;
  LAYER M2 ;
        RECT 4.13 14.14 5.33 14.42 ;
  LAYER M2 ;
        RECT 4.13 8.26 5.33 8.54 ;
  LAYER M2 ;
        RECT 3.7 14.56 4.9 14.84 ;
  LAYER M2 ;
        RECT 3.7 10.36 4.9 10.64 ;
  LAYER M3 ;
        RECT 5.02 8.24 5.3 14.44 ;
  LAYER M1 ;
        RECT 7.185 11.255 7.435 14.785 ;
  LAYER M1 ;
        RECT 7.185 9.995 7.435 11.005 ;
  LAYER M1 ;
        RECT 7.185 7.895 7.435 8.905 ;
  LAYER M1 ;
        RECT 7.615 11.255 7.865 14.785 ;
  LAYER M1 ;
        RECT 6.755 11.255 7.005 14.785 ;
  LAYER M2 ;
        RECT 6.71 14.14 7.91 14.42 ;
  LAYER M2 ;
        RECT 6.71 8.26 7.91 8.54 ;
  LAYER M2 ;
        RECT 7.14 14.56 8.34 14.84 ;
  LAYER M2 ;
        RECT 7.14 10.36 8.34 10.64 ;
  LAYER M3 ;
        RECT 6.74 8.24 7.02 14.44 ;
  END 
END CP

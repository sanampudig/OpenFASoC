MACRO PD
  ORIGIN 0 0 ;
  FOREIGN PD 0 0 ;
  SIZE 23.65 BY 15.12 ;
  PIN 0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 3.3 0.68 3.58 6.88 ;
      LAYER M3 ;
        RECT 1.58 0.68 1.86 6.88 ;
      LAYER M3 ;
        RECT 3.3 3.595 3.58 3.965 ;
      LAYER M2 ;
        RECT 1.72 3.64 3.44 3.92 ;
      LAYER M3 ;
        RECT 1.58 3.595 1.86 3.965 ;
      LAYER M3 ;
        RECT 6.74 0.68 7.02 6.88 ;
      LAYER M3 ;
        RECT 8.46 0.68 8.74 6.88 ;
      LAYER M3 ;
        RECT 6.74 3.595 7.02 3.965 ;
      LAYER M2 ;
        RECT 6.88 3.64 8.6 3.92 ;
      LAYER M3 ;
        RECT 8.46 3.595 8.74 3.965 ;
      LAYER M3 ;
        RECT 16.2 1.1 16.48 6.88 ;
      LAYER M2 ;
        RECT 11.44 0.7 12.64 0.98 ;
      LAYER M3 ;
        RECT 3.3 3.595 3.58 3.965 ;
      LAYER M4 ;
        RECT 3.44 3.38 6.88 4.18 ;
      LAYER M3 ;
        RECT 6.74 3.595 7.02 3.965 ;
      LAYER M3 ;
        RECT 8.46 3.595 8.74 3.965 ;
      LAYER M4 ;
        RECT 8.6 3.38 16.34 4.18 ;
      LAYER M3 ;
        RECT 16.2 3.595 16.48 3.965 ;
      LAYER M4 ;
        RECT 11.875 3.38 12.205 4.18 ;
      LAYER M3 ;
        RECT 11.9 0.84 12.18 3.78 ;
      LAYER M2 ;
        RECT 11.88 0.7 12.2 0.98 ;
    END
  END 0
  PIN 1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 3.3 8.24 3.58 14.44 ;
      LAYER M3 ;
        RECT 1.58 8.24 1.86 14.44 ;
      LAYER M3 ;
        RECT 3.3 11.155 3.58 11.525 ;
      LAYER M2 ;
        RECT 1.72 11.2 3.44 11.48 ;
      LAYER M3 ;
        RECT 1.58 11.155 1.86 11.525 ;
      LAYER M3 ;
        RECT 6.74 8.24 7.02 14.44 ;
      LAYER M3 ;
        RECT 8.46 8.24 8.74 14.44 ;
      LAYER M3 ;
        RECT 6.74 11.155 7.02 11.525 ;
      LAYER M2 ;
        RECT 6.88 11.2 8.6 11.48 ;
      LAYER M3 ;
        RECT 8.46 11.155 8.74 11.525 ;
      LAYER M2 ;
        RECT 18.75 7.84 19.95 8.12 ;
      LAYER M2 ;
        RECT 14.45 7.84 15.65 8.12 ;
      LAYER M3 ;
        RECT 3.3 11.155 3.58 11.525 ;
      LAYER M4 ;
        RECT 3.44 10.94 6.88 11.74 ;
      LAYER M3 ;
        RECT 6.74 11.155 7.02 11.525 ;
      LAYER M3 ;
        RECT 8.46 8.635 8.74 9.005 ;
      LAYER M2 ;
        RECT 8.6 8.68 18.06 8.96 ;
      LAYER M1 ;
        RECT 17.935 7.98 18.185 8.82 ;
      LAYER M2 ;
        RECT 18.06 7.84 18.92 8.12 ;
      LAYER M2 ;
        RECT 14.89 8.68 15.21 8.96 ;
      LAYER M3 ;
        RECT 14.91 7.98 15.19 8.82 ;
      LAYER M2 ;
        RECT 14.89 7.84 15.21 8.12 ;
    END
  END 1
  PIN UP
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 0.26 7 1.46 7.28 ;
      LAYER M2 ;
        RECT 0.26 7.84 1.46 8.12 ;
      LAYER M2 ;
        RECT 0.7 7 1.02 7.28 ;
      LAYER M3 ;
        RECT 0.72 7.14 1 7.98 ;
      LAYER M2 ;
        RECT 0.7 7.84 1.02 8.12 ;
    END
  END UP
  PIN DOWN
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 8.86 7 10.06 7.28 ;
      LAYER M2 ;
        RECT 8.86 7.84 10.06 8.12 ;
      LAYER M2 ;
        RECT 9.3 7 9.62 7.28 ;
      LAYER M3 ;
        RECT 9.32 7.14 9.6 7.98 ;
      LAYER M2 ;
        RECT 9.3 7.84 9.62 8.12 ;
    END
  END DOWN
  PIN CLK2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 17.46 4.48 18.66 4.76 ;
      LAYER M3 ;
        RECT 11.9 7.82 12.18 12.34 ;
      LAYER M2 ;
        RECT 13.16 2.8 14.36 3.08 ;
      LAYER M2 ;
        RECT 14.45 12.04 15.65 12.32 ;
      LAYER M2 ;
        RECT 11.44 2.8 12.64 3.08 ;
      LAYER M2 ;
        RECT 12.04 4.48 17.63 4.76 ;
      LAYER M3 ;
        RECT 11.9 4.62 12.18 7.98 ;
      LAYER M2 ;
        RECT 13.6 4.48 13.92 4.76 ;
      LAYER M3 ;
        RECT 13.62 2.94 13.9 4.62 ;
      LAYER M2 ;
        RECT 13.6 2.8 13.92 3.08 ;
      LAYER M3 ;
        RECT 11.9 11.155 12.18 11.525 ;
      LAYER M2 ;
        RECT 12.04 11.2 12.9 11.48 ;
      LAYER M1 ;
        RECT 12.775 11.34 13.025 12.18 ;
      LAYER M2 ;
        RECT 12.9 12.04 14.62 12.32 ;
      LAYER M2 ;
        RECT 12.47 2.8 13.33 3.08 ;
    END
  END CLK2
  PIN CLK1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 16.6 4.9 17.8 5.18 ;
      LAYER M3 ;
        RECT 22.22 7.82 22.5 12.34 ;
      LAYER M2 ;
        RECT 20.04 2.8 21.24 3.08 ;
      LAYER M2 ;
        RECT 16.17 12.04 17.37 12.32 ;
      LAYER M2 ;
        RECT 18.75 12.04 19.95 12.32 ;
      LAYER M2 ;
        RECT 17.63 4.9 22.36 5.18 ;
      LAYER M3 ;
        RECT 22.22 5.04 22.5 7.98 ;
      LAYER M2 ;
        RECT 20.48 4.9 20.8 5.18 ;
      LAYER M3 ;
        RECT 20.5 2.94 20.78 5.04 ;
      LAYER M2 ;
        RECT 20.48 2.8 20.8 3.08 ;
      LAYER M3 ;
        RECT 22.22 12.18 22.5 12.6 ;
      LAYER M2 ;
        RECT 18.06 12.46 22.36 12.74 ;
      LAYER M1 ;
        RECT 17.935 12.18 18.185 12.6 ;
      LAYER M2 ;
        RECT 17.2 12.04 18.06 12.32 ;
      LAYER M2 ;
        RECT 19.19 12.46 19.51 12.74 ;
      LAYER M1 ;
        RECT 19.225 12.18 19.475 12.6 ;
      LAYER M2 ;
        RECT 19.19 12.04 19.51 12.32 ;
    END
  END CLK1
  OBS 
  LAYER M2 ;
        RECT 3.7 2.8 4.9 3.08 ;
  LAYER M2 ;
        RECT 3.7 12.04 4.9 12.32 ;
  LAYER M2 ;
        RECT 3.71 2.8 4.03 3.08 ;
  LAYER M3 ;
        RECT 3.73 2.94 4.01 12.18 ;
  LAYER M2 ;
        RECT 3.71 12.04 4.03 12.32 ;
  LAYER M3 ;
        RECT 21.79 8.24 22.07 14.44 ;
  LAYER M2 ;
        RECT 16.17 7.84 17.37 8.12 ;
  LAYER M2 ;
        RECT 4.57 12.04 4.89 12.32 ;
  LAYER M1 ;
        RECT 4.605 11.76 4.855 12.18 ;
  LAYER M2 ;
        RECT 4.73 11.62 21.93 11.9 ;
  LAYER M3 ;
        RECT 21.79 11.575 22.07 11.945 ;
  LAYER M2 ;
        RECT 16.61 11.62 16.93 11.9 ;
  LAYER M3 ;
        RECT 16.63 7.98 16.91 11.76 ;
  LAYER M2 ;
        RECT 16.61 7.84 16.93 8.12 ;
  LAYER M1 ;
        RECT 4.605 11.675 4.855 11.845 ;
  LAYER M2 ;
        RECT 4.56 11.62 4.9 11.9 ;
  LAYER M1 ;
        RECT 4.605 12.095 4.855 12.265 ;
  LAYER M2 ;
        RECT 4.56 12.04 4.9 12.32 ;
  LAYER M2 ;
        RECT 21.77 11.62 22.09 11.9 ;
  LAYER M3 ;
        RECT 21.79 11.6 22.07 11.92 ;
  LAYER M1 ;
        RECT 4.605 11.675 4.855 11.845 ;
  LAYER M2 ;
        RECT 4.56 11.62 4.9 11.9 ;
  LAYER M1 ;
        RECT 4.605 12.095 4.855 12.265 ;
  LAYER M2 ;
        RECT 4.56 12.04 4.9 12.32 ;
  LAYER M2 ;
        RECT 21.77 11.62 22.09 11.9 ;
  LAYER M3 ;
        RECT 21.79 11.6 22.07 11.92 ;
  LAYER M1 ;
        RECT 4.605 11.675 4.855 11.845 ;
  LAYER M2 ;
        RECT 4.56 11.62 4.9 11.9 ;
  LAYER M1 ;
        RECT 4.605 12.095 4.855 12.265 ;
  LAYER M2 ;
        RECT 4.56 12.04 4.9 12.32 ;
  LAYER M2 ;
        RECT 16.61 7.84 16.93 8.12 ;
  LAYER M3 ;
        RECT 16.63 7.82 16.91 8.14 ;
  LAYER M2 ;
        RECT 16.61 11.62 16.93 11.9 ;
  LAYER M3 ;
        RECT 16.63 11.6 16.91 11.92 ;
  LAYER M2 ;
        RECT 21.77 11.62 22.09 11.9 ;
  LAYER M3 ;
        RECT 21.79 11.6 22.07 11.92 ;
  LAYER M1 ;
        RECT 4.605 11.675 4.855 11.845 ;
  LAYER M2 ;
        RECT 4.56 11.62 4.9 11.9 ;
  LAYER M1 ;
        RECT 4.605 12.095 4.855 12.265 ;
  LAYER M2 ;
        RECT 4.56 12.04 4.9 12.32 ;
  LAYER M2 ;
        RECT 16.61 7.84 16.93 8.12 ;
  LAYER M3 ;
        RECT 16.63 7.82 16.91 8.14 ;
  LAYER M2 ;
        RECT 16.61 11.62 16.93 11.9 ;
  LAYER M3 ;
        RECT 16.63 11.6 16.91 11.92 ;
  LAYER M2 ;
        RECT 21.77 11.62 22.09 11.9 ;
  LAYER M3 ;
        RECT 21.79 11.6 22.07 11.92 ;
  LAYER M2 ;
        RECT 5.42 2.8 6.62 3.08 ;
  LAYER M2 ;
        RECT 5.42 12.04 6.62 12.32 ;
  LAYER M2 ;
        RECT 5.43 2.8 5.75 3.08 ;
  LAYER M1 ;
        RECT 5.465 2.94 5.715 12.18 ;
  LAYER M2 ;
        RECT 5.43 12.04 5.75 12.32 ;
  LAYER M3 ;
        RECT 12.33 8.24 12.61 14.44 ;
  LAYER M2 ;
        RECT 11.44 7 12.64 7.28 ;
  LAYER M2 ;
        RECT 6.29 12.04 6.61 12.32 ;
  LAYER M3 ;
        RECT 6.31 12.18 6.59 12.6 ;
  LAYER M2 ;
        RECT 6.45 12.46 12.47 12.74 ;
  LAYER M3 ;
        RECT 12.33 12.415 12.61 12.785 ;
  LAYER M3 ;
        RECT 12.33 7.14 12.61 8.4 ;
  LAYER M2 ;
        RECT 12.31 7 12.63 7.28 ;
  LAYER M2 ;
        RECT 6.29 12.04 6.61 12.32 ;
  LAYER M3 ;
        RECT 6.31 12.02 6.59 12.34 ;
  LAYER M2 ;
        RECT 6.29 12.46 6.61 12.74 ;
  LAYER M3 ;
        RECT 6.31 12.44 6.59 12.76 ;
  LAYER M2 ;
        RECT 12.31 12.46 12.63 12.74 ;
  LAYER M3 ;
        RECT 12.33 12.44 12.61 12.76 ;
  LAYER M2 ;
        RECT 6.29 12.04 6.61 12.32 ;
  LAYER M3 ;
        RECT 6.31 12.02 6.59 12.34 ;
  LAYER M2 ;
        RECT 6.29 12.46 6.61 12.74 ;
  LAYER M3 ;
        RECT 6.31 12.44 6.59 12.76 ;
  LAYER M2 ;
        RECT 12.31 12.46 12.63 12.74 ;
  LAYER M3 ;
        RECT 12.33 12.44 12.61 12.76 ;
  LAYER M2 ;
        RECT 6.29 12.04 6.61 12.32 ;
  LAYER M3 ;
        RECT 6.31 12.02 6.59 12.34 ;
  LAYER M2 ;
        RECT 6.29 12.46 6.61 12.74 ;
  LAYER M3 ;
        RECT 6.31 12.44 6.59 12.76 ;
  LAYER M2 ;
        RECT 12.31 7 12.63 7.28 ;
  LAYER M3 ;
        RECT 12.33 6.98 12.61 7.3 ;
  LAYER M2 ;
        RECT 12.31 12.46 12.63 12.74 ;
  LAYER M3 ;
        RECT 12.33 12.44 12.61 12.76 ;
  LAYER M2 ;
        RECT 6.29 12.04 6.61 12.32 ;
  LAYER M3 ;
        RECT 6.31 12.02 6.59 12.34 ;
  LAYER M2 ;
        RECT 6.29 12.46 6.61 12.74 ;
  LAYER M3 ;
        RECT 6.31 12.44 6.59 12.76 ;
  LAYER M2 ;
        RECT 12.31 7 12.63 7.28 ;
  LAYER M3 ;
        RECT 12.33 6.98 12.61 7.3 ;
  LAYER M2 ;
        RECT 12.31 12.46 12.63 12.74 ;
  LAYER M3 ;
        RECT 12.33 12.44 12.61 12.76 ;
  LAYER M2 ;
        RECT 17.46 0.28 18.66 0.56 ;
  LAYER M3 ;
        RECT 19.64 0.68 19.92 6.88 ;
  LAYER M2 ;
        RECT 18.49 0.28 19.78 0.56 ;
  LAYER M3 ;
        RECT 19.64 0.42 19.92 0.84 ;
  LAYER M2 ;
        RECT 19.62 0.28 19.94 0.56 ;
  LAYER M3 ;
        RECT 19.64 0.26 19.92 0.58 ;
  LAYER M2 ;
        RECT 19.62 0.28 19.94 0.56 ;
  LAYER M3 ;
        RECT 19.64 0.26 19.92 0.58 ;
  LAYER M2 ;
        RECT 16.6 0.7 17.8 0.98 ;
  LAYER M3 ;
        RECT 14.48 0.68 14.76 6.88 ;
  LAYER M2 ;
        RECT 15.48 0.7 16.77 0.98 ;
  LAYER M1 ;
        RECT 15.355 0.84 15.605 1.26 ;
  LAYER M2 ;
        RECT 14.62 1.12 15.48 1.4 ;
  LAYER M3 ;
        RECT 14.48 1.075 14.76 1.445 ;
  LAYER M1 ;
        RECT 15.355 0.755 15.605 0.925 ;
  LAYER M2 ;
        RECT 15.31 0.7 15.65 0.98 ;
  LAYER M1 ;
        RECT 15.355 1.175 15.605 1.345 ;
  LAYER M2 ;
        RECT 15.31 1.12 15.65 1.4 ;
  LAYER M2 ;
        RECT 14.46 1.12 14.78 1.4 ;
  LAYER M3 ;
        RECT 14.48 1.1 14.76 1.42 ;
  LAYER M1 ;
        RECT 15.355 0.755 15.605 0.925 ;
  LAYER M2 ;
        RECT 15.31 0.7 15.65 0.98 ;
  LAYER M1 ;
        RECT 15.355 1.175 15.605 1.345 ;
  LAYER M2 ;
        RECT 15.31 1.12 15.65 1.4 ;
  LAYER M2 ;
        RECT 14.46 1.12 14.78 1.4 ;
  LAYER M3 ;
        RECT 14.48 1.1 14.76 1.42 ;
  LAYER M2 ;
        RECT 20.04 7 21.24 7.28 ;
  LAYER M3 ;
        RECT 17.49 8.24 17.77 14.44 ;
  LAYER M3 ;
        RECT 20.07 8.24 20.35 14.44 ;
  LAYER M2 ;
        RECT 17.63 7 20.21 7.28 ;
  LAYER M3 ;
        RECT 17.49 7.14 17.77 8.4 ;
  LAYER M2 ;
        RECT 20.05 7 20.37 7.28 ;
  LAYER M3 ;
        RECT 20.07 7.14 20.35 8.4 ;
  LAYER M2 ;
        RECT 17.47 7 17.79 7.28 ;
  LAYER M3 ;
        RECT 17.49 6.98 17.77 7.3 ;
  LAYER M2 ;
        RECT 17.47 7 17.79 7.28 ;
  LAYER M3 ;
        RECT 17.49 6.98 17.77 7.3 ;
  LAYER M2 ;
        RECT 17.47 7 17.79 7.28 ;
  LAYER M3 ;
        RECT 17.49 6.98 17.77 7.3 ;
  LAYER M2 ;
        RECT 20.05 7 20.37 7.28 ;
  LAYER M3 ;
        RECT 20.07 6.98 20.35 7.3 ;
  LAYER M2 ;
        RECT 17.47 7 17.79 7.28 ;
  LAYER M3 ;
        RECT 17.49 6.98 17.77 7.3 ;
  LAYER M2 ;
        RECT 20.05 7 20.37 7.28 ;
  LAYER M3 ;
        RECT 20.07 6.98 20.35 7.3 ;
  LAYER M2 ;
        RECT 13.16 7 14.36 7.28 ;
  LAYER M3 ;
        RECT 14.05 8.24 14.33 14.44 ;
  LAYER M2 ;
        RECT 11.01 6.58 12.21 6.86 ;
  LAYER M2 ;
        RECT 14.03 7 14.35 7.28 ;
  LAYER M3 ;
        RECT 14.05 7.14 14.33 8.4 ;
  LAYER M2 ;
        RECT 13.17 7 13.49 7.28 ;
  LAYER M1 ;
        RECT 13.205 6.3 13.455 7.14 ;
  LAYER M2 ;
        RECT 12.9 6.16 13.33 6.44 ;
  LAYER M1 ;
        RECT 12.775 6.3 13.025 6.72 ;
  LAYER M2 ;
        RECT 12.04 6.58 12.9 6.86 ;
  LAYER M2 ;
        RECT 14.03 7 14.35 7.28 ;
  LAYER M3 ;
        RECT 14.05 6.98 14.33 7.3 ;
  LAYER M2 ;
        RECT 14.03 7 14.35 7.28 ;
  LAYER M3 ;
        RECT 14.05 6.98 14.33 7.3 ;
  LAYER M1 ;
        RECT 12.775 6.215 13.025 6.385 ;
  LAYER M2 ;
        RECT 12.73 6.16 13.07 6.44 ;
  LAYER M1 ;
        RECT 12.775 6.635 13.025 6.805 ;
  LAYER M2 ;
        RECT 12.73 6.58 13.07 6.86 ;
  LAYER M1 ;
        RECT 13.205 6.215 13.455 6.385 ;
  LAYER M2 ;
        RECT 13.16 6.16 13.5 6.44 ;
  LAYER M1 ;
        RECT 13.205 7.055 13.455 7.225 ;
  LAYER M2 ;
        RECT 13.16 7 13.5 7.28 ;
  LAYER M2 ;
        RECT 14.03 7 14.35 7.28 ;
  LAYER M3 ;
        RECT 14.05 6.98 14.33 7.3 ;
  LAYER M1 ;
        RECT 12.775 6.215 13.025 6.385 ;
  LAYER M2 ;
        RECT 12.73 6.16 13.07 6.44 ;
  LAYER M1 ;
        RECT 12.775 6.635 13.025 6.805 ;
  LAYER M2 ;
        RECT 12.73 6.58 13.07 6.86 ;
  LAYER M1 ;
        RECT 13.205 6.215 13.455 6.385 ;
  LAYER M2 ;
        RECT 13.16 6.16 13.5 6.44 ;
  LAYER M1 ;
        RECT 13.205 7.055 13.455 7.225 ;
  LAYER M2 ;
        RECT 13.16 7 13.5 7.28 ;
  LAYER M2 ;
        RECT 14.03 7 14.35 7.28 ;
  LAYER M3 ;
        RECT 14.05 6.98 14.33 7.3 ;
  LAYER M2 ;
        RECT 3.7 7 4.9 7.28 ;
  LAYER M2 ;
        RECT 3.7 7.84 4.9 8.12 ;
  LAYER M2 ;
        RECT 4.14 7 4.46 7.28 ;
  LAYER M3 ;
        RECT 4.16 7.14 4.44 7.98 ;
  LAYER M2 ;
        RECT 4.14 7.84 4.46 8.12 ;
  LAYER M2 ;
        RECT 0.26 2.8 1.46 3.08 ;
  LAYER M2 ;
        RECT 0.26 12.04 1.46 12.32 ;
  LAYER M2 ;
        RECT 0.27 2.8 0.59 3.08 ;
  LAYER M1 ;
        RECT 0.305 2.94 0.555 12.18 ;
  LAYER M2 ;
        RECT 0.27 12.04 0.59 12.32 ;
  LAYER M3 ;
        RECT 4.16 7.375 4.44 7.745 ;
  LAYER M2 ;
        RECT 0.43 7.42 4.3 7.7 ;
  LAYER M1 ;
        RECT 0.305 7.475 0.555 7.645 ;
  LAYER M1 ;
        RECT 0.305 7.475 0.555 7.645 ;
  LAYER M2 ;
        RECT 0.26 7.42 0.6 7.7 ;
  LAYER M2 ;
        RECT 4.14 7.42 4.46 7.7 ;
  LAYER M3 ;
        RECT 4.16 7.4 4.44 7.72 ;
  LAYER M1 ;
        RECT 0.305 7.475 0.555 7.645 ;
  LAYER M2 ;
        RECT 0.26 7.42 0.6 7.7 ;
  LAYER M2 ;
        RECT 4.14 7.42 4.46 7.7 ;
  LAYER M3 ;
        RECT 4.16 7.4 4.44 7.72 ;
  LAYER M1 ;
        RECT 3.745 3.695 3.995 7.225 ;
  LAYER M1 ;
        RECT 3.745 2.435 3.995 3.445 ;
  LAYER M1 ;
        RECT 3.745 0.335 3.995 1.345 ;
  LAYER M1 ;
        RECT 4.175 3.695 4.425 7.225 ;
  LAYER M1 ;
        RECT 3.315 3.695 3.565 7.225 ;
  LAYER M2 ;
        RECT 3.27 0.7 4.47 0.98 ;
  LAYER M2 ;
        RECT 3.27 6.58 4.47 6.86 ;
  LAYER M2 ;
        RECT 3.7 7 4.9 7.28 ;
  LAYER M2 ;
        RECT 3.7 2.8 4.9 3.08 ;
  LAYER M3 ;
        RECT 3.3 0.68 3.58 6.88 ;
  LAYER M1 ;
        RECT 3.745 7.895 3.995 11.425 ;
  LAYER M1 ;
        RECT 3.745 11.675 3.995 12.685 ;
  LAYER M1 ;
        RECT 3.745 13.775 3.995 14.785 ;
  LAYER M1 ;
        RECT 4.175 7.895 4.425 11.425 ;
  LAYER M1 ;
        RECT 3.315 7.895 3.565 11.425 ;
  LAYER M2 ;
        RECT 3.27 14.14 4.47 14.42 ;
  LAYER M2 ;
        RECT 3.27 8.26 4.47 8.54 ;
  LAYER M2 ;
        RECT 3.7 7.84 4.9 8.12 ;
  LAYER M2 ;
        RECT 3.7 12.04 4.9 12.32 ;
  LAYER M3 ;
        RECT 3.3 8.24 3.58 14.44 ;
  LAYER M1 ;
        RECT 1.165 3.695 1.415 7.225 ;
  LAYER M1 ;
        RECT 1.165 2.435 1.415 3.445 ;
  LAYER M1 ;
        RECT 1.165 0.335 1.415 1.345 ;
  LAYER M1 ;
        RECT 0.735 3.695 0.985 7.225 ;
  LAYER M1 ;
        RECT 1.595 3.695 1.845 7.225 ;
  LAYER M2 ;
        RECT 0.69 0.7 1.89 0.98 ;
  LAYER M2 ;
        RECT 0.69 6.58 1.89 6.86 ;
  LAYER M2 ;
        RECT 0.26 7 1.46 7.28 ;
  LAYER M2 ;
        RECT 0.26 2.8 1.46 3.08 ;
  LAYER M3 ;
        RECT 1.58 0.68 1.86 6.88 ;
  LAYER M1 ;
        RECT 1.165 7.895 1.415 11.425 ;
  LAYER M1 ;
        RECT 1.165 11.675 1.415 12.685 ;
  LAYER M1 ;
        RECT 1.165 13.775 1.415 14.785 ;
  LAYER M1 ;
        RECT 0.735 7.895 0.985 11.425 ;
  LAYER M1 ;
        RECT 1.595 7.895 1.845 11.425 ;
  LAYER M2 ;
        RECT 0.69 14.14 1.89 14.42 ;
  LAYER M2 ;
        RECT 0.69 8.26 1.89 8.54 ;
  LAYER M2 ;
        RECT 0.26 7.84 1.46 8.12 ;
  LAYER M2 ;
        RECT 0.26 12.04 1.46 12.32 ;
  LAYER M3 ;
        RECT 1.58 8.24 1.86 14.44 ;
  LAYER M2 ;
        RECT 5.42 7 6.62 7.28 ;
  LAYER M2 ;
        RECT 5.42 7.84 6.62 8.12 ;
  LAYER M2 ;
        RECT 5.86 7 6.18 7.28 ;
  LAYER M3 ;
        RECT 5.88 7.14 6.16 7.98 ;
  LAYER M2 ;
        RECT 5.86 7.84 6.18 8.12 ;
  LAYER M2 ;
        RECT 8.86 2.8 10.06 3.08 ;
  LAYER M2 ;
        RECT 8.86 12.04 10.06 12.32 ;
  LAYER M2 ;
        RECT 8.87 2.8 9.19 3.08 ;
  LAYER M3 ;
        RECT 8.89 2.94 9.17 12.18 ;
  LAYER M2 ;
        RECT 8.87 12.04 9.19 12.32 ;
  LAYER M3 ;
        RECT 5.88 7.375 6.16 7.745 ;
  LAYER M2 ;
        RECT 6.02 7.42 9.03 7.7 ;
  LAYER M3 ;
        RECT 8.89 7.375 9.17 7.745 ;
  LAYER M2 ;
        RECT 5.86 7.42 6.18 7.7 ;
  LAYER M3 ;
        RECT 5.88 7.4 6.16 7.72 ;
  LAYER M2 ;
        RECT 8.87 7.42 9.19 7.7 ;
  LAYER M3 ;
        RECT 8.89 7.4 9.17 7.72 ;
  LAYER M2 ;
        RECT 5.86 7.42 6.18 7.7 ;
  LAYER M3 ;
        RECT 5.88 7.4 6.16 7.72 ;
  LAYER M2 ;
        RECT 8.87 7.42 9.19 7.7 ;
  LAYER M3 ;
        RECT 8.89 7.4 9.17 7.72 ;
  LAYER M1 ;
        RECT 6.325 3.695 6.575 7.225 ;
  LAYER M1 ;
        RECT 6.325 2.435 6.575 3.445 ;
  LAYER M1 ;
        RECT 6.325 0.335 6.575 1.345 ;
  LAYER M1 ;
        RECT 5.895 3.695 6.145 7.225 ;
  LAYER M1 ;
        RECT 6.755 3.695 7.005 7.225 ;
  LAYER M2 ;
        RECT 5.85 0.7 7.05 0.98 ;
  LAYER M2 ;
        RECT 5.85 6.58 7.05 6.86 ;
  LAYER M2 ;
        RECT 5.42 7 6.62 7.28 ;
  LAYER M2 ;
        RECT 5.42 2.8 6.62 3.08 ;
  LAYER M3 ;
        RECT 6.74 0.68 7.02 6.88 ;
  LAYER M1 ;
        RECT 6.325 7.895 6.575 11.425 ;
  LAYER M1 ;
        RECT 6.325 11.675 6.575 12.685 ;
  LAYER M1 ;
        RECT 6.325 13.775 6.575 14.785 ;
  LAYER M1 ;
        RECT 5.895 7.895 6.145 11.425 ;
  LAYER M1 ;
        RECT 6.755 7.895 7.005 11.425 ;
  LAYER M2 ;
        RECT 5.85 14.14 7.05 14.42 ;
  LAYER M2 ;
        RECT 5.85 8.26 7.05 8.54 ;
  LAYER M2 ;
        RECT 5.42 7.84 6.62 8.12 ;
  LAYER M2 ;
        RECT 5.42 12.04 6.62 12.32 ;
  LAYER M3 ;
        RECT 6.74 8.24 7.02 14.44 ;
  LAYER M1 ;
        RECT 8.905 3.695 9.155 7.225 ;
  LAYER M1 ;
        RECT 8.905 2.435 9.155 3.445 ;
  LAYER M1 ;
        RECT 8.905 0.335 9.155 1.345 ;
  LAYER M1 ;
        RECT 9.335 3.695 9.585 7.225 ;
  LAYER M1 ;
        RECT 8.475 3.695 8.725 7.225 ;
  LAYER M2 ;
        RECT 8.43 0.7 9.63 0.98 ;
  LAYER M2 ;
        RECT 8.43 6.58 9.63 6.86 ;
  LAYER M2 ;
        RECT 8.86 7 10.06 7.28 ;
  LAYER M2 ;
        RECT 8.86 2.8 10.06 3.08 ;
  LAYER M3 ;
        RECT 8.46 0.68 8.74 6.88 ;
  LAYER M1 ;
        RECT 8.905 7.895 9.155 11.425 ;
  LAYER M1 ;
        RECT 8.905 11.675 9.155 12.685 ;
  LAYER M1 ;
        RECT 8.905 13.775 9.155 14.785 ;
  LAYER M1 ;
        RECT 9.335 7.895 9.585 11.425 ;
  LAYER M1 ;
        RECT 8.475 7.895 8.725 11.425 ;
  LAYER M2 ;
        RECT 8.43 14.14 9.63 14.42 ;
  LAYER M2 ;
        RECT 8.43 8.26 9.63 8.54 ;
  LAYER M2 ;
        RECT 8.86 7.84 10.06 8.12 ;
  LAYER M2 ;
        RECT 8.86 12.04 10.06 12.32 ;
  LAYER M3 ;
        RECT 8.46 8.24 8.74 14.44 ;
  LAYER M1 ;
        RECT 17.505 0.335 17.755 3.865 ;
  LAYER M1 ;
        RECT 17.505 4.115 17.755 5.125 ;
  LAYER M1 ;
        RECT 17.505 6.215 17.755 7.225 ;
  LAYER M1 ;
        RECT 17.935 0.335 18.185 3.865 ;
  LAYER M1 ;
        RECT 17.075 0.335 17.325 3.865 ;
  LAYER M1 ;
        RECT 16.645 0.335 16.895 3.865 ;
  LAYER M1 ;
        RECT 16.645 4.115 16.895 5.125 ;
  LAYER M1 ;
        RECT 16.645 6.215 16.895 7.225 ;
  LAYER M1 ;
        RECT 16.215 0.335 16.465 3.865 ;
  LAYER M2 ;
        RECT 16.17 6.58 17.8 6.86 ;
  LAYER M2 ;
        RECT 16.17 1.12 18.23 1.4 ;
  LAYER M2 ;
        RECT 17.46 0.28 18.66 0.56 ;
  LAYER M2 ;
        RECT 16.6 0.7 17.8 0.98 ;
  LAYER M2 ;
        RECT 17.46 4.48 18.66 4.76 ;
  LAYER M2 ;
        RECT 16.6 4.9 17.8 5.18 ;
  LAYER M3 ;
        RECT 16.2 1.1 16.48 6.88 ;
  LAYER M1 ;
        RECT 11.915 7.895 12.165 11.425 ;
  LAYER M1 ;
        RECT 11.915 11.675 12.165 12.685 ;
  LAYER M1 ;
        RECT 11.915 13.775 12.165 14.785 ;
  LAYER M1 ;
        RECT 11.485 7.895 11.735 11.425 ;
  LAYER M1 ;
        RECT 12.345 7.895 12.595 11.425 ;
  LAYER M2 ;
        RECT 11.01 12.04 12.21 12.32 ;
  LAYER M2 ;
        RECT 11.01 7.84 12.21 8.12 ;
  LAYER M2 ;
        RECT 11.44 14.14 12.64 14.42 ;
  LAYER M2 ;
        RECT 11.44 8.26 12.64 8.54 ;
  LAYER M3 ;
        RECT 11.9 7.82 12.18 12.34 ;
  LAYER M3 ;
        RECT 12.33 8.24 12.61 14.44 ;
  LAYER M1 ;
        RECT 22.235 7.895 22.485 11.425 ;
  LAYER M1 ;
        RECT 22.235 11.675 22.485 12.685 ;
  LAYER M1 ;
        RECT 22.235 13.775 22.485 14.785 ;
  LAYER M1 ;
        RECT 22.665 7.895 22.915 11.425 ;
  LAYER M1 ;
        RECT 21.805 7.895 22.055 11.425 ;
  LAYER M2 ;
        RECT 22.19 12.04 23.39 12.32 ;
  LAYER M2 ;
        RECT 22.19 7.84 23.39 8.12 ;
  LAYER M2 ;
        RECT 21.76 14.14 22.96 14.42 ;
  LAYER M2 ;
        RECT 21.76 8.26 22.96 8.54 ;
  LAYER M3 ;
        RECT 22.22 7.82 22.5 12.34 ;
  LAYER M3 ;
        RECT 21.79 8.24 22.07 14.44 ;
  LAYER M1 ;
        RECT 20.085 3.695 20.335 7.225 ;
  LAYER M1 ;
        RECT 20.085 2.435 20.335 3.445 ;
  LAYER M1 ;
        RECT 20.085 0.335 20.335 1.345 ;
  LAYER M1 ;
        RECT 20.515 3.695 20.765 7.225 ;
  LAYER M1 ;
        RECT 19.655 3.695 19.905 7.225 ;
  LAYER M2 ;
        RECT 19.61 0.7 20.81 0.98 ;
  LAYER M2 ;
        RECT 19.61 6.58 20.81 6.86 ;
  LAYER M2 ;
        RECT 20.04 7 21.24 7.28 ;
  LAYER M2 ;
        RECT 20.04 2.8 21.24 3.08 ;
  LAYER M3 ;
        RECT 19.64 0.68 19.92 6.88 ;
  LAYER M1 ;
        RECT 14.065 3.695 14.315 7.225 ;
  LAYER M1 ;
        RECT 14.065 2.435 14.315 3.445 ;
  LAYER M1 ;
        RECT 14.065 0.335 14.315 1.345 ;
  LAYER M1 ;
        RECT 13.635 3.695 13.885 7.225 ;
  LAYER M1 ;
        RECT 14.495 3.695 14.745 7.225 ;
  LAYER M2 ;
        RECT 13.59 0.7 14.79 0.98 ;
  LAYER M2 ;
        RECT 13.59 6.58 14.79 6.86 ;
  LAYER M2 ;
        RECT 13.16 7 14.36 7.28 ;
  LAYER M2 ;
        RECT 13.16 2.8 14.36 3.08 ;
  LAYER M3 ;
        RECT 14.48 0.68 14.76 6.88 ;
  LAYER M1 ;
        RECT 17.075 7.895 17.325 11.425 ;
  LAYER M1 ;
        RECT 17.075 11.675 17.325 12.685 ;
  LAYER M1 ;
        RECT 17.075 13.775 17.325 14.785 ;
  LAYER M1 ;
        RECT 16.645 7.895 16.895 11.425 ;
  LAYER M1 ;
        RECT 17.505 7.895 17.755 11.425 ;
  LAYER M2 ;
        RECT 16.6 14.14 17.8 14.42 ;
  LAYER M2 ;
        RECT 16.6 8.26 17.8 8.54 ;
  LAYER M2 ;
        RECT 16.17 7.84 17.37 8.12 ;
  LAYER M2 ;
        RECT 16.17 12.04 17.37 12.32 ;
  LAYER M3 ;
        RECT 17.49 8.24 17.77 14.44 ;
  LAYER M1 ;
        RECT 19.655 7.895 19.905 11.425 ;
  LAYER M1 ;
        RECT 19.655 11.675 19.905 12.685 ;
  LAYER M1 ;
        RECT 19.655 13.775 19.905 14.785 ;
  LAYER M1 ;
        RECT 19.225 7.895 19.475 11.425 ;
  LAYER M1 ;
        RECT 20.085 7.895 20.335 11.425 ;
  LAYER M2 ;
        RECT 19.18 14.14 20.38 14.42 ;
  LAYER M2 ;
        RECT 19.18 8.26 20.38 8.54 ;
  LAYER M2 ;
        RECT 18.75 7.84 19.95 8.12 ;
  LAYER M2 ;
        RECT 18.75 12.04 19.95 12.32 ;
  LAYER M3 ;
        RECT 20.07 8.24 20.35 14.44 ;
  LAYER M1 ;
        RECT 14.495 7.895 14.745 11.425 ;
  LAYER M1 ;
        RECT 14.495 11.675 14.745 12.685 ;
  LAYER M1 ;
        RECT 14.495 13.775 14.745 14.785 ;
  LAYER M1 ;
        RECT 14.925 7.895 15.175 11.425 ;
  LAYER M1 ;
        RECT 14.065 7.895 14.315 11.425 ;
  LAYER M2 ;
        RECT 14.02 14.14 15.22 14.42 ;
  LAYER M2 ;
        RECT 14.02 8.26 15.22 8.54 ;
  LAYER M2 ;
        RECT 14.45 7.84 15.65 8.12 ;
  LAYER M2 ;
        RECT 14.45 12.04 15.65 12.32 ;
  LAYER M3 ;
        RECT 14.05 8.24 14.33 14.44 ;
  LAYER M1 ;
        RECT 11.485 3.695 11.735 7.225 ;
  LAYER M1 ;
        RECT 11.485 2.435 11.735 3.445 ;
  LAYER M1 ;
        RECT 11.485 0.335 11.735 1.345 ;
  LAYER M1 ;
        RECT 11.915 3.695 12.165 7.225 ;
  LAYER M1 ;
        RECT 11.055 3.695 11.305 7.225 ;
  LAYER M2 ;
        RECT 11.44 0.7 12.64 0.98 ;
  LAYER M2 ;
        RECT 11.44 7 12.64 7.28 ;
  LAYER M2 ;
        RECT 11.44 2.8 12.64 3.08 ;
  LAYER M2 ;
        RECT 11.01 6.58 12.21 6.86 ;
  END 
END PD
